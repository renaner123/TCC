pll_2M_inst : pll_2M PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
